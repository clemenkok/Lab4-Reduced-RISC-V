module name #(
    parameters
) (
    port_list
);
    
endmodule